module decoder (
  input logic [3:0] binary,

  output logic [15:0] one_hot
);
  always_comb begin 
    one_hot = 16'b0000_0000_0000_0000;
      case (binary)
      4'b0000: one_hot = 16'b0000_0000_0000_0001; // 0
      4'b0001: one_hot = 16'b0000_0000_0000_0010; // 1
      4'b0010: one_hot = 16'b0000_0000_0000_0100; // 2
      4'b0011: one_hot = 16'b0000_0000_0000_1000; // 3
      4'b0100: one_hot = 16'b0000_0000_0001_0000; // 4
      4'b0101: one_hot = 16'b0000_0000_0010_0000; // 5
      4'b0110: one_hot = 16'b0000_0000_0100_0000; // 6
      4'b0111: one_hot = 16'b0000_0000_1000_0000; // 7
      4'b1000: one_hot = 16'b0000_0001_0000_0000; // 8
      4'b1001: one_hot = 16'b0000_0010_0000_0000; // 9
      4'b1010: one_hot = 16'b0000_0100_0000_0000; // 10
      4'b1011: one_hot = 16'b0000_1000_0000_0000; // 11
      4'b1100: one_hot = 16'b0001_0000_0000_0000; // 12
      4'b1101: one_hot = 16'b0010_0000_0000_0000; // 13
      4'b1110: one_hot = 16'b0100_0000_0000_0000; // 14
      4'b1111: one_hot = 16'b1000_0000_0000_0000; // 15
      default: one_hot = 16'b0000_0000_0000_0000; // other conditions
    endcase  
  end

endmodule