module decoder (
  input logic [3:0] binary,

  output logic [15:0] one_hot
);

  //add description here 
  //

endmodule