module decoder (
  input logic [3:0] binary,

  output logic [15:0] one_hot
);

  // description here 111


endmodule

module decoder (
  input logic [3:0] binary,

  output logic [15:0] one_hot
);

  // description here 111

endmodule